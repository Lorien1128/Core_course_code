`timescale 1ns / 1ps
`define IDLE 2'b00
`define LOAD 2'b01
`define CNT  2'b10
`define INT  2'b11

`define ctrl   mem[0]
`define preset mem[1]
`define count  mem[2]
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:43:39 12/28/2017 
// Design Name: 
// Module Name:    TC 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module TC(
    input clk,
    input reset,
    input [31:2] Addr,
    input WE,
    input [31:0] Din,
    output [31:0] Dout,
    output IRQ	//����ж�����
    );

	reg [1:0] state;
	reg [31:0] mem [2:0];	//mem[0]:CTRL, mem[1]:PRESET, mem[2]:COUNT
	
	reg _IRQ;
	assign IRQ = `ctrl[3] & _IRQ;	//ctrl[3]==1���������ж�
	
	assign Dout = mem[Addr[3:2]];	//Addr��[3:2]λ��ʾҪ��д�ļĴ������
	
	wire [31:0] load = Addr[3:2] == 0 ? {28'h0, Din[3:0]} : Din;	//дCTRL�Ĵ���ʱֻд����λ
	
	integer i;
	always @(posedge clk) begin
		if(reset) begin		//��λΪ0
			state <= 0; 
			for(i = 0; i < 3; i = i+1) mem[i] <= 0;
			_IRQ <= 0;
		end
		else if(WE) begin
			// $display("%d@: *%h <= %h", $time, {Addr, 2'b00}, load);
			mem[Addr[3:2]] <= load;	//д�Ĵ���
		end
		else begin
			case(state)
				`IDLE : if(`ctrl[0]) begin	//����̬��������ʹ����Чʱ��������̬�������ж�
					state <= `LOAD;
					_IRQ <= 1'b0;
				end
				`LOAD : begin		//����̬������������Ϊ��ʼֵ���������̬
					`count <= `preset;
					state <= `CNT;
				end
				`CNT  : 			//����̬
					if(`ctrl[0]) begin	//������ʹ����Чʱ��countÿ������-1
						if(`count > 1) `count <= `count-1;
						else begin	//count����0ʱ�����ж�̬
							`count <= 0;
							state <= `INT;
							_IRQ <= 1'b1;
						end
					end
					else state <= `IDLE;	//������ʹ����Чʱ�ص�����̬
				default : begin		//`INT���ж�̬
					if(`ctrl[2:1] == 2'b00) `ctrl[0] <= 1'b0;	//ģʽ0��������ʹ����0�������ж�ֱ��ʹ�ܱ���1
					else _IRQ <= 1'b0;			//ģʽ1��ֱ��ֹͣ�ж�
					state <= `IDLE;			//����ģʽ���ص�����̬
				end
			endcase
		end
	end

endmodule
